// Defines for BlackIce-II
