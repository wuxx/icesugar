// Defines for iCEBreaker
`define SPI_FLASH
`define INTERNAL_OSC
