// Defines for ECP5 evaluation board
